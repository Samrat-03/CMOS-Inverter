magic
tech sky130A
timestamp 1709920053
<< nwell >>
rect -300 0 0 415
<< nmos >>
rect -155 -200 -140 -100
<< pmos >>
rect -155 50 -140 250
<< ndiff >>
rect -200 -110 -155 -100
rect -200 -190 -190 -110
rect -170 -190 -155 -110
rect -200 -200 -155 -190
rect -140 -110 -95 -100
rect -140 -190 -125 -110
rect -105 -190 -95 -110
rect -140 -200 -95 -190
<< pdiff >>
rect -200 240 -155 250
rect -200 60 -190 240
rect -170 60 -155 240
rect -200 50 -155 60
rect -140 240 -95 250
rect -140 60 -125 240
rect -105 60 -95 240
rect -140 50 -95 60
<< ndiffc >>
rect -190 -190 -170 -110
rect -125 -190 -105 -110
<< pdiffc >>
rect -190 60 -170 240
rect -125 60 -105 240
<< psubdiff >>
rect -220 -245 -70 -230
rect -220 -270 -205 -245
rect -85 -270 -70 -245
rect -220 -285 -70 -270
<< nsubdiff >>
rect -225 375 -75 390
rect -225 350 -210 375
rect -90 350 -75 375
rect -225 335 -75 350
<< psubdiffcont >>
rect -205 -270 -85 -245
<< nsubdiffcont >>
rect -210 350 -90 375
<< poly >>
rect -155 250 -140 305
rect -155 -15 -140 50
rect -190 -25 -140 -15
rect -190 -45 -185 -25
rect -165 -45 -140 -25
rect -190 -55 -140 -45
rect -155 -100 -140 -55
rect -155 -215 -140 -200
<< polycont >>
rect -185 -45 -165 -25
<< locali >>
rect -225 380 -75 390
rect -225 375 -185 380
rect -125 375 -75 380
rect -225 350 -210 375
rect -90 350 -75 375
rect -225 345 -185 350
rect -125 345 -75 350
rect -225 335 -75 345
rect -200 240 -160 335
rect -200 60 -190 240
rect -170 60 -160 240
rect -200 50 -160 60
rect -135 240 -95 250
rect -135 60 -125 240
rect -105 60 -95 240
rect -190 -25 -155 -15
rect -190 -45 -185 -25
rect -165 -45 -155 -25
rect -190 -55 -155 -45
rect -135 -25 -95 60
rect -135 -45 -125 -25
rect -105 -45 -95 -25
rect -200 -110 -160 -100
rect -200 -190 -190 -110
rect -170 -190 -160 -110
rect -200 -230 -160 -190
rect -135 -110 -95 -45
rect -135 -190 -125 -110
rect -105 -190 -95 -110
rect -135 -200 -95 -190
rect -220 -240 -70 -230
rect -220 -245 -185 -240
rect -125 -245 -70 -240
rect -220 -270 -205 -245
rect -85 -270 -70 -245
rect -220 -275 -185 -270
rect -125 -275 -70 -270
rect -220 -285 -70 -275
<< viali >>
rect -185 375 -125 380
rect -185 350 -125 375
rect -185 345 -125 350
rect -185 -45 -165 -25
rect -125 -45 -105 -25
rect -185 -245 -125 -240
rect -185 -270 -125 -245
rect -185 -275 -125 -270
<< metal1 >>
rect -455 380 170 390
rect -455 345 -185 380
rect -125 345 170 380
rect -455 335 170 345
rect -430 -25 -155 -15
rect -430 -45 -185 -25
rect -165 -45 -155 -25
rect -430 -55 -155 -45
rect -135 -25 120 -15
rect -135 -45 -125 -25
rect -105 -45 120 -25
rect -135 -55 120 -45
rect -455 -240 170 -230
rect -455 -275 -185 -240
rect -125 -275 170 -240
rect -455 -285 170 -275
<< labels >>
rlabel metal1 95 360 95 360 1 vcc
rlabel metal1 55 -260 55 -260 1 gnd
rlabel metal1 -115 -55 120 -15 1 vout
rlabel metal1 -310 -40 -310 -40 1 vin
<< end >>
